module fsm(input clk);



endmodule