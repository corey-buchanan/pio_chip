module pio_core(
    input clk,
    input rst,
    input [31:0] gpio_input,
    output reg [31:0] core_output,
    output reg [31:0] core_drive
    );

    reg [4:0] pc;
    reg [15:0] instruction;
    reg [15:0] data_in;
    reg [4:0] write_addr;
    reg write_en;

    // Remove when spi is wired up
    initial begin
        write_addr = 5'b00000;
        write_en = 0;
    end

    // Add the other FSMs later
    fsm fsm(
        .clk(clk),
        .rst(rst),
        .instruction(instruction),
        .pc(pc)
        // TODO - add fifo push/pop en, status, etc.
    );

    // TODO - Wire these up to the FSMs
    reg [31:0] fsm_output [3:0];
    reg [31:0] fsm_drive [3:0];

    // TODO - Wire signals up to fsm
    // These FIFOs are reversable, will need to store direction
    // the names right now refer to their default direction
    // I'll have a look at the docs to see if that's the best way
    // to name these fifos
    reg [31:0] tx_data_in;
    reg tx_push_en;
    reg tx_pop_en;
    reg [31:0] tx_data_out;
    reg [1:0] tx_status;
    reg [2:0] tx_fifo_count;

    reg [31:0] rx_data_in;
    reg rx_push_en;
    reg rx_pop_en;
    reg [31:0] rx_data_out;
    reg [1:0] rx_status;
    reg [2:0] rx_fifo_count;

    fifo tx_fifo (
        .clk(clk),
        .rst(rst),
        .data_in(tx_data_in),
        .push_en(tx_push_en),
        .pop_en(tx_pop_en),
        .data_out(tx_data_out),
        .status(tx_status),
        .fifo_count(tx_fifo_count)
    );

    fifo rx_fifo (
        .clk(clk),
        .rst(rst),
        .data_in(gpio_input),
        .push_en(1),
        .pop_en(1),
        .data_out(rx_data_out),
        .status(rx_status),
        .fifo_count(rx_fifo_count)
    );

    // TODO Add OSR

    fsm_output_arbitrator fsm_output_arbitrator(
        .fsm_output(fsm_output),
        .fsm_drive(fsm_drive),
        .core_output(core_output),
        .core_drive(core_drive)
    );

    instruction_regfile instruction_regfile(
        .clk(clk),
        .rst(rst),
        .data_in(data_in),
        .write_addr(write_addr),
        .write_en(write_en),
        .read_addr(pc),
        .data_out(instruction)
    );

endmodule